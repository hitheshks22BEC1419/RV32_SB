
//module pipeline3 #(parameter WIDTH = 32)(
//    input wire[WIDTH-1:0] a,b,
//    input wire add_sub, //1:sub
    
//)